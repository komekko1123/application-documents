module Shifter(in, shamt, out);
	input [31:0] in ; 
	input [4:0] shamt ; //  8 = 3, 16 = 4, 32 = 5 
	output [31:0] out ;
	wire [31:0] x,y,z,w;
	// 16 bit shift right
	Mux_2to1  s4_31 (.in0(in[31]),.in1(1'b0),.sel(shamt[4]),.out(w[31]) );
	Mux_2to1  s4_30 (.in0(in[30]),.in1(1'b0),.sel(shamt[4]),.out(w[30]) );
	Mux_2to1  s4_29 (.in0(in[29]),.in1(1'b0),.sel(shamt[4]),.out(w[29]) );
	Mux_2to1  s4_28 (.in0(in[28]),.in1(1'b0),.sel(shamt[4]),.out(w[28]) );
	Mux_2to1  s4_27 (.in0(in[27]),.in1(1'b0),.sel(shamt[4]),.out(w[27]) );
	Mux_2to1  s4_26 (.in0(in[26]),.in1(1'b0),.sel(shamt[4]),.out(w[26]) );
	Mux_2to1  s4_25 (.in0(in[25]),.in1(1'b0),.sel(shamt[4]),.out(w[25]) );
	Mux_2to1  s4_24 (.in0(in[24]),.in1(1'b0),.sel(shamt[4]),.out(w[24]) );
	Mux_2to1  s4_23 (.in0(in[23]),.in1(1'b0),.sel(shamt[4]),.out(w[23]) );
	Mux_2to1  s4_22 (.in0(in[22]),.in1(1'b0),.sel(shamt[4]),.out(w[22]) );
	Mux_2to1  s4_21 (.in0(in[21]),.in1(1'b0),.sel(shamt[4]),.out(w[21]) );
	Mux_2to1  s4_20 (.in0(in[20]),.in1(1'b0),.sel(shamt[4]),.out(w[20]) );
	Mux_2to1  s4_19 (.in0(in[19]),.in1(1'b0),.sel(shamt[4]),.out(w[19]) );
	Mux_2to1  s4_18 (.in0(in[18]),.in1(1'b0),.sel(shamt[4]),.out(w[18]) );
	Mux_2to1  s4_17 (.in0(in[17]),.in1(1'b0),.sel(shamt[4]),.out(w[17]) );
	Mux_2to1  s4_16 (.in0(in[16]),.in1(1'b0),.sel(shamt[4]),.out(w[16]) );
	Mux_2to1  s4_15 (.in0(in[15]),.in1(in[31]),.sel(shamt[4]),.out(w[15]) );
	Mux_2to1  s4_14 (.in0(in[14]),.in1(in[30]),.sel(shamt[4]),.out(w[14]) );
	Mux_2to1  s4_13 (.in0(in[13]),.in1(in[29]),.sel(shamt[4]),.out(w[13]) );
	Mux_2to1  s4_12 (.in0(in[12]),.in1(in[28]),.sel(shamt[4]),.out(w[12]) );
	Mux_2to1  s4_11 (.in0(in[11]),.in1(in[27]),.sel(shamt[4]),.out(w[11]) );
	Mux_2to1  s4_10 (.in0(in[10]),.in1(in[26]),.sel(shamt[4]),.out(w[10]) );
	Mux_2to1  s4_9 (.in0(in[9]),.in1(in[25]),.sel(shamt[4]),.out(w[9]) );
	Mux_2to1  s4_8 (.in0(in[8]),.in1(in[24]),.sel(shamt[4]),.out(w[8]) );
	Mux_2to1  s4_7 (.in0(in[7]),.in1(in[23]),.sel(shamt[4]),.out(w[7]) );
	Mux_2to1  s4_6 (.in0(in[6]),.in1(in[22]),.sel(shamt[4]),.out(w[6]) );
	Mux_2to1  s4_5 (.in0(in[5]),.in1(in[21]),.sel(shamt[4]),.out(w[5]) );
	Mux_2to1  s4_4 (.in0(in[4]),.in1(in[20]),.sel(shamt[4]),.out(w[4]) );
	Mux_2to1  s4_3 (.in0(in[3]),.in1(in[19]),.sel(shamt[4]),.out(w[3]) );
	Mux_2to1  s4_2 (.in0(in[2]),.in1(in[18]),.sel(shamt[4]),.out(w[2]) );
	Mux_2to1  s4_1 (.in0(in[1]),.in1(in[17]),.sel(shamt[4]),.out(w[1]) );
	Mux_2to1  s4_0 (.in0(in[0]),.in1(in[16]),.sel(shamt[4]),.out(w[0]) );
	
	// 8 bit shift right
	Mux_2to1  s3_31 (.in0(w[31]),.in1(1'b0),.sel(shamt[3]),.out(z[31]) );
	Mux_2to1  s3_30 (.in0(w[30]),.in1(1'b0),.sel(shamt[3]),.out(z[30]) );
	Mux_2to1  s3_29 (.in0(w[29]),.in1(1'b0),.sel(shamt[3]),.out(z[29]) );
	Mux_2to1  s3_28 (.in0(w[28]),.in1(1'b0),.sel(shamt[3]),.out(z[28]) );
	Mux_2to1  s3_27 (.in0(w[27]),.in1(1'b0),.sel(shamt[3]),.out(z[27]) );
	Mux_2to1  s3_26 (.in0(w[26]),.in1(1'b0),.sel(shamt[3]),.out(z[26]) );
	Mux_2to1  s3_25 (.in0(w[25]),.in1(1'b0),.sel(shamt[3]),.out(z[25]) );
	Mux_2to1  s3_24 (.in0(w[24]),.in1(1'b0),.sel(shamt[3]),.out(z[24]) );
	Mux_2to1  s3_23 (.in0(w[23]),.in1(w[31]),.sel(shamt[3]),.out(z[23]) );
	Mux_2to1  s3_22 (.in0(w[22]),.in1(w[30]),.sel(shamt[3]),.out(z[22]) );
	Mux_2to1  s3_21 (.in0(w[21]),.in1(w[29]),.sel(shamt[3]),.out(z[21]) );
	Mux_2to1  s3_20 (.in0(w[20]),.in1(w[28]),.sel(shamt[3]),.out(z[20]) );
	Mux_2to1  s3_19 (.in0(w[19]),.in1(w[27]),.sel(shamt[3]),.out(z[19]) );
	Mux_2to1  s3_18 (.in0(w[18]),.in1(w[26]),.sel(shamt[3]),.out(z[18]) );
	Mux_2to1  s3_17 (.in0(w[17]),.in1(w[25]),.sel(shamt[3]),.out(z[17]) );
	Mux_2to1  s3_16 (.in0(w[16]),.in1(w[24]),.sel(shamt[3]),.out(z[16]) );
	Mux_2to1  s3_15 (.in0(w[15]),.in1(w[23]),.sel(shamt[3]),.out(z[15]) );
	Mux_2to1  s3_14 (.in0(w[14]),.in1(w[22]),.sel(shamt[3]),.out(z[14]) );
	Mux_2to1  s3_13 (.in0(w[13]),.in1(w[21]),.sel(shamt[3]),.out(z[13]) );
	Mux_2to1  s3_12 (.in0(w[12]),.in1(w[20]),.sel(shamt[3]),.out(z[12]) );
	Mux_2to1  s3_11 (.in0(w[11]),.in1(w[19]),.sel(shamt[3]),.out(z[11]) );
	Mux_2to1  s3_10 (.in0(w[10]),.in1(w[18]),.sel(shamt[3]),.out(z[10]) );
	Mux_2to1  s3_9 (.in0(w[9]),.in1(w[17]),.sel(shamt[3]),.out(z[9]) );
	Mux_2to1  s3_8 (.in0(w[8]),.in1(w[16]),.sel(shamt[3]),.out(z[8]) );
	Mux_2to1  s3_7 (.in0(w[7]),.in1(w[15]),.sel(shamt[3]),.out(z[7]) );
	Mux_2to1  s3_6 (.in0(w[6]),.in1(w[14]),.sel(shamt[3]),.out(z[6]) );
	Mux_2to1  s3_5 (.in0(w[5]),.in1(w[13]),.sel(shamt[3]),.out(z[5]) );
	Mux_2to1  s3_4 (.in0(w[4]),.in1(w[12]),.sel(shamt[3]),.out(z[4]) );
	Mux_2to1  s3_3 (.in0(w[3]),.in1(w[11]),.sel(shamt[3]),.out(z[3]) );
	Mux_2to1  s3_2 (.in0(w[2]),.in1(w[10]),.sel(shamt[3]),.out(z[2]) );
	Mux_2to1  s3_1 (.in0(w[1]),.in1(w[9]),.sel(shamt[3]),.out(z[1]) );
	Mux_2to1  s3_0 (.in0(w[0]),.in1(w[8]),.sel(shamt[3]),.out(z[0]) );
	
	// 4 bit shift right
	Mux_2to1  s2_31 (.in0(z[31]),.in1(1'b0),.sel(shamt[2]),.out(y[31]) );
	Mux_2to1  s2_30 (.in0(z[30]),.in1(1'b0),.sel(shamt[2]),.out(y[30]) );
	Mux_2to1  s2_29 (.in0(z[29]),.in1(1'b0),.sel(shamt[2]),.out(y[29]) );
	Mux_2to1  s2_28 (.in0(z[28]),.in1(1'b0),.sel(shamt[2]),.out(y[28]) );
	Mux_2to1  s2_27 (.in0(z[27]),.in1(z[31]),.sel(shamt[2]),.out(y[27]) );
	Mux_2to1  s2_26 (.in0(z[26]),.in1(z[30]),.sel(shamt[2]),.out(y[26]) );
	Mux_2to1  s2_25 (.in0(z[25]),.in1(z[29]),.sel(shamt[2]),.out(y[25]) );
	Mux_2to1  s2_24 (.in0(z[24]),.in1(z[28]),.sel(shamt[2]),.out(y[24]) );
	Mux_2to1  s2_23 (.in0(z[23]),.in1(z[27]),.sel(shamt[2]),.out(y[23]) );
	Mux_2to1  s2_22 (.in0(z[22]),.in1(z[26]),.sel(shamt[2]),.out(y[22]) );
	Mux_2to1  s2_21 (.in0(z[21]),.in1(z[25]),.sel(shamt[2]),.out(y[21]) );
	Mux_2to1  s2_20 (.in0(z[20]),.in1(z[24]),.sel(shamt[2]),.out(y[20]) );
	Mux_2to1  s2_19 (.in0(z[19]),.in1(z[23]),.sel(shamt[2]),.out(y[19]) );
	Mux_2to1  s2_18 (.in0(z[18]),.in1(z[22]),.sel(shamt[2]),.out(y[18]) );
	Mux_2to1  s2_17 (.in0(z[17]),.in1(z[21]),.sel(shamt[2]),.out(y[17]) );
	Mux_2to1  s2_16 (.in0(z[16]),.in1(z[20]),.sel(shamt[2]),.out(y[16]) );
	Mux_2to1  s2_15 (.in0(z[15]),.in1(z[19]),.sel(shamt[2]),.out(y[15]) );
	Mux_2to1  s2_14 (.in0(z[14]),.in1(z[18]),.sel(shamt[2]),.out(y[14]) );
	Mux_2to1  s2_13 (.in0(z[13]),.in1(z[17]),.sel(shamt[2]),.out(y[13]) );
	Mux_2to1  s2_12 (.in0(z[12]),.in1(z[16]),.sel(shamt[2]),.out(y[12]) );
	Mux_2to1  s2_11 (.in0(z[11]),.in1(z[15]),.sel(shamt[2]),.out(y[11]) );
	Mux_2to1  s2_10 (.in0(z[10]),.in1(z[14]),.sel(shamt[2]),.out(y[10]) );
	Mux_2to1  s2_9 (.in0(z[9]),.in1(z[13]),.sel(shamt[2]),.out(y[9]) );
	Mux_2to1  s2_8 (.in0(z[8]),.in1(z[12]),.sel(shamt[2]),.out(y[8]) );
	Mux_2to1  s2_7 (.in0(z[7]),.in1(z[11]),.sel(shamt[2]),.out(y[7]) );
	Mux_2to1  s2_6 (.in0(z[6]),.in1(z[10]),.sel(shamt[2]),.out(y[6]) );
	Mux_2to1  s2_5 (.in0(z[5]),.in1(z[9]),.sel(shamt[2]),.out(y[5]) );
	Mux_2to1  s2_4 (.in0(z[4]),.in1(z[8]),.sel(shamt[2]),.out(y[4]) );
	Mux_2to1  s2_3 (.in0(z[3]),.in1(z[7]),.sel(shamt[2]),.out(y[3]) );
	Mux_2to1  s2_2 (.in0(z[2]),.in1(z[6]),.sel(shamt[2]),.out(y[2]) );
	Mux_2to1  s2_1 (.in0(z[1]),.in1(z[5]),.sel(shamt[2]),.out(y[1]) );
	Mux_2to1  s2_0 (.in0(z[0]),.in1(z[4]),.sel(shamt[2]),.out(y[0]) );

	//2 bit shift right

	Mux_2to1  s1_31 (.in0(y[31]),.in1(1'b0),.sel(shamt[1]),.out(x[31]) );
	Mux_2to1  s1_30 (.in0(y[30]),.in1(1'b0),.sel(shamt[1]),.out(x[30]) );
	Mux_2to1  s1_29 (.in0(y[29]),.in1(y[31]),.sel(shamt[1]),.out(x[29]) );
	Mux_2to1  s1_28 (.in0(y[28]),.in1(y[30]),.sel(shamt[1]),.out(x[28]) );
	Mux_2to1  s1_27 (.in0(y[27]),.in1(y[29]),.sel(shamt[1]),.out(x[27]) );
	Mux_2to1  s1_26 (.in0(y[26]),.in1(y[28]),.sel(shamt[1]),.out(x[26]) );
	Mux_2to1  s1_25 (.in0(y[25]),.in1(y[27]),.sel(shamt[1]),.out(x[25]) );
	Mux_2to1  s1_24 (.in0(y[24]),.in1(y[26]),.sel(shamt[1]),.out(x[24]) );
	Mux_2to1  s1_23 (.in0(y[23]),.in1(y[25]),.sel(shamt[1]),.out(x[23]) );
	Mux_2to1  s1_22 (.in0(y[22]),.in1(y[24]),.sel(shamt[1]),.out(x[22]) );
	Mux_2to1  s1_21 (.in0(y[21]),.in1(y[23]),.sel(shamt[1]),.out(x[21]) );
	Mux_2to1  s1_20 (.in0(y[20]),.in1(y[22]),.sel(shamt[1]),.out(x[20]) );
	Mux_2to1  s1_19 (.in0(y[19]),.in1(y[21]),.sel(shamt[1]),.out(x[19]) );
	Mux_2to1  s1_18 (.in0(y[18]),.in1(y[20]),.sel(shamt[1]),.out(x[18]) );
	Mux_2to1  s1_17 (.in0(y[17]),.in1(y[19]),.sel(shamt[1]),.out(x[17]) );
	Mux_2to1  s1_16 (.in0(y[16]),.in1(y[18]),.sel(shamt[1]),.out(x[16]) );
	Mux_2to1  s1_15 (.in0(y[15]),.in1(y[17]),.sel(shamt[1]),.out(x[15]) );
	Mux_2to1  s1_14 (.in0(y[14]),.in1(y[16]),.sel(shamt[1]),.out(x[14]) );
	Mux_2to1  s1_13 (.in0(y[13]),.in1(y[15]),.sel(shamt[1]),.out(x[13]) );
	Mux_2to1  s1_12 (.in0(y[12]),.in1(y[14]),.sel(shamt[1]),.out(x[12]) );
	Mux_2to1  s1_11 (.in0(y[11]),.in1(y[13]),.sel(shamt[1]),.out(x[11]) );
	Mux_2to1  s1_10 (.in0(y[10]),.in1(y[12]),.sel(shamt[1]),.out(x[10]) );
	Mux_2to1  s1_9 (.in0(y[9]),.in1(y[11]),.sel(shamt[1]),.out(x[9]) );
	Mux_2to1  s1_8 (.in0(y[8]),.in1(y[10]),.sel(shamt[1]),.out(x[8]) );
	Mux_2to1  s1_7 (.in0(y[7]),.in1(y[9]),.sel(shamt[1]),.out(x[7]) );
	Mux_2to1  s1_6 (.in0(y[6]),.in1(y[8]),.sel(shamt[1]),.out(x[6]) );
	Mux_2to1  s1_5 (.in0(y[5]),.in1(y[7]),.sel(shamt[1]),.out(x[5]) );
	Mux_2to1  s1_4 (.in0(y[4]),.in1(y[6]),.sel(shamt[1]),.out(x[4]) );
	Mux_2to1  s1_3 (.in0(y[3]),.in1(y[5]),.sel(shamt[1]),.out(x[3]) );
	Mux_2to1  s1_2 (.in0(y[2]),.in1(y[4]),.sel(shamt[1]),.out(x[2]) );
	Mux_2to1  s1_1 (.in0(y[1]),.in1(y[3]),.sel(shamt[1]),.out(x[1]) );
	Mux_2to1  s1_0 (.in0(y[0]),.in1(y[2]),.sel(shamt[1]),.out(x[0]) );	


	//1 bit shift right
	Mux_2to1  s0_31 (.in0(x[31]),.in1(1'b0),.sel(shamt[0]),.out(out[31]) );
	Mux_2to1  s0_30 (.in0(x[30]),.in1(x[31]),.sel(shamt[0]),.out(out[30]) );
	Mux_2to1  s0_29 (.in0(x[29]),.in1(x[30]),.sel(shamt[0]),.out(out[29]) );
	Mux_2to1  s0_28 (.in0(x[28]),.in1(x[29]),.sel(shamt[0]),.out(out[28]) );
	Mux_2to1  s0_27 (.in0(x[27]),.in1(x[28]),.sel(shamt[0]),.out(out[27]) );
	Mux_2to1  s0_26 (.in0(x[26]),.in1(x[27]),.sel(shamt[0]),.out(out[26]) );
	Mux_2to1  s0_25 (.in0(x[25]),.in1(x[26]),.sel(shamt[0]),.out(out[25]) );
	Mux_2to1  s0_24 (.in0(x[24]),.in1(x[25]),.sel(shamt[0]),.out(out[24]) );
	Mux_2to1  s0_23 (.in0(x[23]),.in1(x[24]),.sel(shamt[0]),.out(out[23]) );
	Mux_2to1  s0_22 (.in0(x[22]),.in1(x[23]),.sel(shamt[0]),.out(out[22]) );
	Mux_2to1  s0_21 (.in0(x[21]),.in1(x[22]),.sel(shamt[0]),.out(out[21]) );
	Mux_2to1  s0_20 (.in0(x[20]),.in1(x[21]),.sel(shamt[0]),.out(out[20]) );
	Mux_2to1  s0_19 (.in0(x[19]),.in1(x[20]),.sel(shamt[0]),.out(out[19]) );
	Mux_2to1  s0_18 (.in0(x[18]),.in1(x[19]),.sel(shamt[0]),.out(out[18]) );
	Mux_2to1  s0_17 (.in0(x[17]),.in1(x[18]),.sel(shamt[0]),.out(out[17]) );
	Mux_2to1  s0_16 (.in0(x[16]),.in1(x[17]),.sel(shamt[0]),.out(out[16]) );
	Mux_2to1  s0_15 (.in0(x[15]),.in1(x[16]),.sel(shamt[0]),.out(out[15]) );
	Mux_2to1  s0_14 (.in0(x[14]),.in1(x[15]),.sel(shamt[0]),.out(out[14]) );
	Mux_2to1  s0_13 (.in0(x[13]),.in1(x[14]),.sel(shamt[0]),.out(out[13]) );
	Mux_2to1  s0_12 (.in0(x[12]),.in1(x[13]),.sel(shamt[0]),.out(out[12]) );
	Mux_2to1  s0_11 (.in0(x[11]),.in1(x[12]),.sel(shamt[0]),.out(out[11]) );
	Mux_2to1  s0_10 (.in0(x[10]),.in1(x[11]),.sel(shamt[0]),.out(out[10]) );
	Mux_2to1  s0_9 (.in0(x[9]),.in1(x[10]),.sel(shamt[0]),.out(out[9]) );
	Mux_2to1  s0_8 (.in0(x[8]),.in1(x[9]),.sel(shamt[0]),.out(out[8]) );
	Mux_2to1  s0_7 (.in0(x[7]),.in1(x[8]),.sel(shamt[0]),.out(out[7]) );
	Mux_2to1  s0_6 (.in0(x[6]),.in1(x[7]),.sel(shamt[0]),.out(out[6]) );
	Mux_2to1  s0_5 (.in0(x[5]),.in1(x[6]),.sel(shamt[0]),.out(out[5]) );
	Mux_2to1  s0_4 (.in0(x[4]),.in1(x[5]),.sel(shamt[0]),.out(out[4]) );
	Mux_2to1  s0_3 (.in0(x[3]),.in1(x[4]),.sel(shamt[0]),.out(out[3]) );
	Mux_2to1  s0_2 (.in0(x[2]),.in1(x[3]),.sel(shamt[0]),.out(out[2]) );
	Mux_2to1  s0_1 (.in0(x[1]),.in1(x[2]),.sel(shamt[0]),.out(out[1]) );
	Mux_2to1  s0_0 (.in0(x[0]),.in1(x[1]),.sel(shamt[0]),.out(out[0]) );

endmodule
